`timescale 1ps/1ns


module register_logic (
    input clk,
    input enable,
    input [4:0] Data,
    output reg [4:0] Q
);
    // Module implementation goes here
endmodule
