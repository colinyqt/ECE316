`timescale 1ps/1ns

module full_adder (
    input A, B, Cin,
    output S, Cout
);
    // Module implementation goes here
endmodule


module RCA_4bits (
    input clk,
    input enable,
    input [3:0] A, B,
    input Cin,
    output [4:0] Q
);
    // Module implementation goes here
endmodule